--	Package File Template
--
--	Purpose: This package defines supplemental types, subtypes, 
--		 constants, and functions 


library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_arith.ALL;

package modules is

  
  type t_muxN is array(natural range <>) of std_logic_vector(7 downto 0);
 
end modules;


package body modules is

end modules;
